module Half_Adder(input in1,input in2,output sum, output carry);

 carry=in1&in2;
 sum=in1^in2;
 
 endmodule 